
`ifndef BUS_SVH
`define BUS_SVH


`include "bus_trans.sv"

`include "bus_source_agent.sv"
`include "bus_source_seq_lib.sv"
`include "bus_destination_agent.sv"

`endif //  `ifndef BUS_SVH

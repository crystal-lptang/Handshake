
`ifndef BUS_PKG_SV
`define BUS_PKG_SV

package bus_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "bus.svh"

endpackage : bus_pkg

   
`endif //  `ifndef BUS_PKG_SV
